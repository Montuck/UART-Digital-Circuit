`timescale 1ns / 1ps
`default_nettype none
/***************************************************************************
*
* Module: FourFunctions
*
* Author: Trevor Wiseman
* Class: ECEN 220, Section 2, Fall 2021
* Date: 09/22/21
*
* Description: LAB 3 Structural SV
*
*
****************************************************************************/

module FourFunctions(

    );
endmodule
